library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sumador_completo is
    Port ( a,b,cin : in  STD_LOGIC;
           s,cout : out  STD_LOGIC);
end sumador_completo;

architecture Behavioral of sumador_completo is

begin


end Behavioral;

